library IEEE;
use IEEE.std_logic_1164.all;
use ieee.numeric_std.all;

entity memoriaROM is
   generic (
          dataWidth: natural := 13;
          addrWidth: natural := 8
    );
   port (
          Endereco : in std_logic_vector (addrWidth-1 DOWNTO 0);
          Dado : out std_logic_vector (dataWidth-1 DOWNTO 0)
    );
end entity;

architecture assincrona of memoriaROM is

  type blocoMemoria is array(0 TO 2**addrWidth - 1) of std_logic_vector(dataWidth-1 DOWNTO 0);
  
  constant NOP  : std_logic_vector(3 downto 0) := "0000";
  constant LDA  : std_logic_vector(3 downto 0) := "0001";
  constant SOMA : std_logic_vector(3 downto 0) := "0010";
  constant SUB  : std_logic_vector(3 downto 0) := "0011";
  constant LDI : std_logic_vector(3 downto 0) := "0100";
  constant STA : std_logic_vector(3 downto 0) := "0101";
  constant JMP : std_logic_vector(3 downto 0) := "0110";
  constant JGE : std_logic_vector(3 downto 0) := "0111";
  constant JEQ : std_logic_vector(3 downto 0) := "1000";
  constant CEQ : std_logic_vector(3 downto 0) := "1001";
  constant JSR : std_logic_vector(3 downto 0) := "1010";
  constant RET : std_logic_vector(3 downto 0) := "1011";
  constant AND1 : std_logic_vector(3 downto 0) := "1100";
  constant JLE : std_logic_vector(3 downto 0) := "1101";
  constant JL : std_logic_vector(3 downto 0) := "1110";
  constant JG : std_logic_vector(3 downto 0) := "1111";

  function initMemory
        return blocoMemoria is variable tmp : blocoMemoria := (others => (others => '0'));
  begin
tmp(0) := LDI & "00" & '0' & x"00";	-- LDI $0 	#Carrega o acumulador com  valor 0
tmp(1) := JSR & "00" & '1' & x"09";	-- JSR @265	#Limpa o display
tmp(2) := JSR & "00" & '1' & x"11";	-- JSR @273	#Limpa os LEDs
tmp(3) := LDI & "00" & '0' & x"00";	-- LDI $0 	#Carrega o acumulador com  valor 0
tmp(4) := STA & "00" & '0' & x"0B";	-- STA @11 	#Zera o valor das unidades
tmp(5) := LDI & "00" & '0' & x"05";	-- LDI $5 
tmp(6) := STA & "00" & '0' & x"0C";	-- STA @12 	#Zera o valor das dezenas
tmp(7) := LDI & "00" & '0' & x"09";	-- LDI $9
tmp(8) := STA & "00" & '0' & x"0D";	-- STA @13 	#Zera o valor das centenas
tmp(9) := LDI & "00" & '0' & x"05";	-- LDI $5
tmp(10) := STA & "00" & '0' & x"0E";	-- STA @14 	#Zera o valor das unidades de milhar
tmp(11) := LDI & "00" & '0' & x"03";	-- LDI $3
tmp(12) := STA & "00" & '0' & x"0F";	-- STA @15 	#Zera o valor das dezenas de milhar
tmp(13) := LDI & "00" & '0' & x"02";	-- LDI $2
tmp(14) := STA & "00" & '0' & x"10";	-- STA @16 	#Zera o valor das centenas de milhar
tmp(15) := LDI & "00" & '0' & x"00";	-- LDI $0 	#Carrega o acumulador com  valor 0
tmp(16) := STA & "00" & '0' & x"11";	-- STA @17 	#Zera a flag de inibir contagem
tmp(17) := STA & "00" & '1' & x"FF";	-- STA @KEY0 	#Limpa a leitura de KEY0
tmp(18) := STA & "00" & '1' & x"FE";	-- STA @KEY1 	#Limpa a leitura de KEY1
tmp(19) := STA & "00" & '1' & x"FD";	-- STA @KEY2 	#Limpa a leitura de KEY2
tmp(20) := STA & "00" & '1' & x"FC";	-- STA @FPGA_RESET 	#Limpa a leitura de FPGA_RESET
tmp(21) := STA & "00" & '0' & x"00";	-- STA @0 	#Criando a constante 0
tmp(22) := LDI & "00" & '0' & x"01";	-- LDI $1 	#Carrega o acumulador com  valor 1
tmp(23) := STA & "00" & '0' & x"01";	-- STA @1 	#Criando a constante 1
tmp(24) := LDI & "00" & '0' & x"02";	-- LDI $2 	#Carrega o acumulador com  valor 2
tmp(25) := STA & "00" & '0' & x"02";	-- STA @2 	#Criando a constante 2
tmp(26) := LDI & "00" & '0' & x"04";	-- LDI $4 	#Carrega o acumulador com  valor 4
tmp(27) := STA & "00" & '0' & x"04";	-- STA @4 	#Criando a constante 4
tmp(28) := LDI & "00" & '0' & x"0F";	-- LDI $15
tmp(29) := STA & "00" & '0' & x"2D";	-- STA @45
tmp(30) := LDI & "00" & '0' & x"05";	-- LDI $5 	#Carrega o acumulador com  valor 5
tmp(31) := STA & "00" & '0' & x"05";	-- STA @5 	#Criando a constante 5
tmp(32) := LDI & "00" & '0' & x"06";	-- LDI $6 	#Carrega o acumulador com  valor 6
tmp(33) := STA & "00" & '0' & x"06";	-- STA @6 	#Criando a constante 6
tmp(34) := LDI & "00" & '0' & x"09";	-- LDI $9 	#Carrega o acumulador com  valor 9
tmp(35) := STA & "00" & '0' & x"09";	-- STA @9 	#Criando a constante 9
tmp(36) := LDI & "00" & '0' & x"0A";	-- LDI $10 	#Carrega o acumulador com  valor 10
tmp(37) := STA & "00" & '0' & x"0A";	-- STA @10 	#Criando a constante 10
tmp(38) := LDI & "00" & '0' & x"00";	-- LDI $0 	#Carrega o acumulador com  valor 0
tmp(39) := STA & "00" & '0' & x"15";	-- STA @21 	#Maximo valor das unidades do limite
tmp(40) := STA & "00" & '0' & x"16";	-- STA @22 	#Maximo valor das dezenas do limite
tmp(41) := STA & "00" & '0' & x"17";	-- STA @23 	#Maximo valor das centenas do limite
tmp(42) := STA & "00" & '0' & x"18";	-- STA @24 	#Maximo valor das unidades de milhar do limite
tmp(43) := STA & "00" & '0' & x"19";	-- STA @25 	#Maximo valor das dezenas de milhar do limite
tmp(44) := LDI & "00" & '0' & x"0A";	-- LDI $10 	#Carrega o acumulador com  valor 10
tmp(45) := STA & "00" & '0' & x"1A";	-- STA @26 	#Maximo valor das centenas de milhar do limite
tmp(46) := LDA & "00" & '1' & x"60";	-- LDA @352 	#Lê KEY0
tmp(47) := AND1 & "00" & '0' & x"01";	-- AND1 @1 	#Mask
tmp(48) := CEQ & "00" & '0' & x"00";	-- CEQ @0 	#Verifica se KEY0 não foi pressionado
tmp(49) := JEQ & "00" & '0' & x"33";	-- JEQ @51	#Se não foi, pula a chamada da subrotina de incremento
tmp(50) := JSR & "00" & '0' & x"45";	-- JSR @69	#Chama a subrotina de incremento
tmp(51) := LDA & "00" & '1' & x"62";	-- LDA @354 	#Lê KEY2
tmp(52) := AND1 & "00" & '0' & x"01";	-- AND1 @1 	#Mask
tmp(53) := CEQ & "00" & '0' & x"00";	-- CEQ @0 	#Verifica se KEY2 não foi pressionado
tmp(54) := JEQ & "00" & '0' & x"38";	-- JEQ @56	#Se não foi, pula a chamada da subrotina de decremento
tmp(55) := JSR & "00" & '0' & x"85";	-- JSR @133	#Chama a subrotina de decremento
tmp(56) := JSR & "00" & '0' & x"C6";	-- JSR @198	#Atualiza o display
tmp(57) := LDA & "00" & '1' & x"61";	-- LDA @353 	#Lê KEY1
tmp(58) := AND1 & "00" & '0' & x"01";	-- AND1 @1 	#Mask
tmp(59) := CEQ & "00" & '0' & x"00";	-- CEQ @0 	#Verifica se KEY1 não foi pressionado
tmp(60) := JEQ & "00" & '0' & x"3E";	-- JEQ @62	#Se não foi, pula a chamada da subrotina de configuracao do limite
tmp(61) := JSR & "00" & '0' & x"D3";	-- JSR @211	#Chama a subrotina de configuracao do limite
tmp(62) := JSR & "00" & '0' & x"E1";	-- JSR @225	#Verifica se o limite foi atingido
tmp(63) := LDA & "00" & '1' & x"64";	-- LDA @356 	#Lê FPGA_RESET
tmp(64) := AND1 & "00" & '0' & x"01";	-- AND1 @1 	#Mask
tmp(65) := CEQ & "00" & '0' & x"00";	-- CEQ @0 	#Verifica se FPGA_RESET não foi pressionado
tmp(66) := JEQ & "00" & '0' & x"44";	-- JEQ @68	#Se não foi, pula a chamada da subrotina de reiniciar contagem
tmp(67) := JSR & "00" & '0' & x"FD";	-- JSR @253	#Chama a subrotina de reiniciar contagem
tmp(68) := JMP & "00" & '0' & x"2E";	-- JMP @46	#Retorna ao inicio do loop
tmp(69) := STA & "00" & '1' & x"FF";	-- STA @KEY0 	#Limpa a leitura de KEY0
tmp(70) := LDA & "00" & '0' & x"11";	-- LDA @17 	#Lê a flag de inibir contagem
tmp(71) := CEQ & "00" & '0' & x"00";	-- CEQ @0 	#Verifica se a contagem não está inibida
tmp(72) := JEQ & "00" & '0' & x"4A";	-- JEQ @74	#Se não estiver, continua a contagem
tmp(73) := RET & "00" & '0' & x"00";	-- RET 	#Se estiver inibida, retorna ao loop principal
tmp(74) := LDI & "00" & '0' & x"01";	-- LDI $1 	#Carrega o acumulador com  valor 1
tmp(75) := SOMA & "00" & '0' & x"0B";	-- SOMA @11 	#Soma o valor das unidades dos segundos com 1
tmp(76) := CEQ & "00" & '0' & x"0A";	-- CEQ @10 	#Verifica se o valor das unidades dos segundos é igual a 10
tmp(77) := JEQ & "00" & '0' & x"50";	-- JEQ @80	#Se sim, incremente a dezena
tmp(78) := STA & "00" & '0' & x"0B";	-- STA @11 	#Armazena o valor das unidades dos segundos
tmp(79) := RET & "00" & '0' & x"00";	-- RET 	#Retorna ao loop principal
tmp(80) := LDI & "00" & '0' & x"00";	-- LDI $0 	#Carrega o acumulador com  valor 0
tmp(81) := STA & "00" & '0' & x"0B";	-- STA @11 	#Zera o valor das unidades dos segundos
tmp(82) := LDI & "00" & '0' & x"01";	-- LDI $1 	#Carrega o acumulador com  valor 1
tmp(83) := SOMA & "00" & '0' & x"0C";	-- SOMA @12 	#Soma o valor das dezenas dos segundos com 1
tmp(84) := CEQ & "00" & '0' & x"06";	-- CEQ @6 	#Verifica se o valor das dezenas dos segundos é igual a 6
tmp(85) := JEQ & "00" & '0' & x"58";	-- JEQ @88	#Se sim, incremente a unidades dos minutos
tmp(86) := STA & "00" & '0' & x"0C";	-- STA @12 	#Armazena o valor das dezenas dos segundos
tmp(87) := RET & "00" & '0' & x"00";	-- RET 	#Retorna ao loop principal
tmp(88) := LDI & "00" & '0' & x"00";	-- LDI $0 	#Carrega o acumulador com  valor 0
tmp(89) := STA & "00" & '0' & x"0C";	-- STA @12 	#Zera o valor das dezenas dos segundos
tmp(90) := LDI & "00" & '0' & x"01";	-- LDI $1 	#Carrega o acumulador com  valor 1
tmp(91) := SOMA & "00" & '0' & x"0D";	-- SOMA @13 	#Soma o valor das unidades dos minutos com 1
tmp(92) := CEQ & "00" & '0' & x"0A";	-- CEQ @10 	#Verifica se o valor das unidades dos minutos é igual a 10
tmp(93) := JEQ & "00" & '0' & x"60";	-- JEQ @96	#Se sim, incremente as dezenas dos minutos
tmp(94) := STA & "00" & '0' & x"0D";	-- STA @13 	#Armazena o valor das unidades dos minutos
tmp(95) := RET & "00" & '0' & x"00";	-- RET 	#Retorna ao loop principal
tmp(96) := LDI & "00" & '0' & x"00";	-- LDI $0 	#Carrega o acumulador com  valor 0
tmp(97) := STA & "00" & '0' & x"0D";	-- STA @13 	#Zera o valor das unidades dos minutos
tmp(98) := LDI & "00" & '0' & x"01";	-- LDI $1 	#Carrega o acumulador com  valor 1
tmp(99) := SOMA & "00" & '0' & x"0E";	-- SOMA @14 	#Soma o valor das dezenas dos minutos com 1
tmp(100) := CEQ & "00" & '0' & x"06";	-- CEQ @6 	#Verifica se o valor das dezenas dos minutos é igual a 6
tmp(101) := JEQ & "00" & '0' & x"68";	-- JEQ @104	#Se sim, incremente as unidades das horas
tmp(102) := STA & "00" & '0' & x"0E";	-- STA @14 	#Armazena o valor das unidades de milhar
tmp(103) := RET & "00" & '0' & x"00";	-- RET 	#Retorna ao loop principal
tmp(104) := LDI & "00" & '0' & x"00";	-- LDI $0 	#Carrega o acumulador com  valor 0
tmp(105) := STA & "00" & '0' & x"0E";	-- STA @14 	#Zera o valor das dezenas dos minutos
tmp(106) := LDI & "00" & '0' & x"01";	-- LDI $1 	#Carrega o acumulador com  valor 1
tmp(107) := SOMA & "00" & '0' & x"0F";	-- SOMA @15 	#Soma o valor das unidades das horas com 1
tmp(108) := CEQ & "00" & '0' & x"0A";	-- CEQ @10 	#Verifica se o valor das unidades das horas é igual a 10
tmp(109) := JEQ & "00" & '0' & x"72";	-- JEQ @114	#Se sim, incremente as unidades das horas
tmp(110) := CEQ & "00" & '0' & x"04";	-- CEQ @4 	#Verifica se o valor das unidades das horas é igual a 4
tmp(111) := JEQ & "00" & '0' & x"78";	-- JEQ @120	#Se sim, cheque se o valor das dezenas de horas é igual a 2
tmp(112) := STA & "00" & '0' & x"0F";	-- STA @15 	#Armazena o valor das unidades das horas
tmp(113) := RET & "00" & '0' & x"00";	-- RET 	#Retorna ao loop principal
tmp(114) := LDI & "00" & '0' & x"00";	-- LDI $0 	#Carrega o acumulador com  valor 0
tmp(115) := STA & "00" & '0' & x"0F";	-- STA @15 	#Zera o valor das unidades das horas
tmp(116) := LDI & "00" & '0' & x"01";	-- LDI $1 	#Carrega o acumulador com  valor 1
tmp(117) := SOMA & "00" & '0' & x"10";	-- SOMA @16 	#Soma o valor das dezenas das horas com 1
tmp(118) := STA & "00" & '0' & x"10";	-- STA @16 	#Armazena o valor das dezenas das horas
tmp(119) := RET & "00" & '0' & x"00";	-- RET 	#Retorna ao loop principal
tmp(120) := LDA & "01" & '0' & x"10";	-- LDA R1, 16 	#Carrega o registrador 1 com o valor das dezenas de horas
tmp(121) := CEQ & "01" & '0' & x"02";	-- CEQ R1, 2 	#Verifica se o valor das dezenas de horas é igual a 2
tmp(122) := JEQ & "00" & '0' & x"7D";	-- JEQ @125	#Se sim, reinicie a contagem
tmp(123) := STA & "00" & '0' & x"0F";	-- STA R0, 15 	#Armazena o valor das unidades de horas
tmp(124) := RET & "00" & '0' & x"00";	-- RET 	#Retorna ao loop principal
tmp(125) := LDI & "00" & '0' & x"00";	-- LDI $0 	#Carrega o acumulador com  valor 0
tmp(126) := STA & "00" & '0' & x"0B";	-- STA @11 	#Armazena o valor das unidades
tmp(127) := STA & "00" & '0' & x"0C";	-- STA @12 	#Armazena o valor das dezenas
tmp(128) := STA & "00" & '0' & x"0D";	-- STA @13 	#Armazena o valor das centenas
tmp(129) := STA & "00" & '0' & x"0E";	-- STA @14 	#Armazena o valor das unidades de milhar
tmp(130) := STA & "00" & '0' & x"0F";	-- STA @15 	#Armazena o valor das dezenas de milhar
tmp(131) := STA & "00" & '0' & x"10";	-- STA @16 	#Armazena o valor das centenas de milhar
tmp(132) := RET & "00" & '0' & x"00";	-- RET 	#Retorna ao loop principal
tmp(133) := STA & "00" & '1' & x"FD";	-- STA @KEY2 	#Limpa a leitura de KEY2
tmp(134) := LDI & "00" & '0' & x"00";	-- LDI $0 	#Carrega o acumulador com  valor 0
tmp(135) := STA & "00" & '0' & x"11";	-- STA @17 	#Zera a flag de inibir contagem
tmp(136) := STA & "00" & '1' & x"01";	-- STA @257 	#Apaga o LED de limite atingido
tmp(137) := STA & "00" & '1' & x"02";	-- STA @258 	#Apaga o LED de overflow
tmp(138) := LDA & "00" & '0' & x"0B";	-- LDA @11 	#Lê o valor das unidades
tmp(139) := CEQ & "00" & '0' & x"00";	-- CEQ @0 	#Verifica se o valor das unidades é igual a 0
tmp(140) := JEQ & "00" & '0' & x"91";	-- JEQ @145	#Se sim, decremente a dezena
tmp(141) := LDA & "00" & '0' & x"0B";	-- LDA @11 	#Carrega o acumulador com  valor 1
tmp(142) := SUB & "00" & '0' & x"01";	-- SUB @1 	#Subtrai 1 do valor das unidades
tmp(143) := STA & "00" & '0' & x"0B";	-- STA @11 	#Armazena o valor das unidades
tmp(144) := RET & "00" & '0' & x"00";	-- RET 	#Retorna ao loop principal
tmp(145) := LDI & "00" & '0' & x"09";	-- LDI $9 	#Carrega o acumulador com  valor 9
tmp(146) := STA & "00" & '0' & x"0B";	-- STA @11 	#Armazena o valor das unidades
tmp(147) := LDA & "00" & '0' & x"0C";	-- LDA @12 	#Lê o valor das dezenas
tmp(148) := CEQ & "00" & '0' & x"00";	-- CEQ @0 	#Verifica se o valor das dezenas é igual a 0
tmp(149) := JEQ & "00" & '0' & x"9A";	-- JEQ @154	#Se sim, decremente a centena
tmp(150) := LDA & "00" & '0' & x"0C";	-- LDA @12 	#Carrega o acumulador com  valor 1
tmp(151) := SUB & "00" & '0' & x"01";	-- SUB @1 	#Subtrai o valor das dezenas com 1
tmp(152) := STA & "00" & '0' & x"0C";	-- STA @12 	#Armazena o valor das dezenas
tmp(153) := RET & "00" & '0' & x"00";	-- RET 	#Retorna ao loop principal
tmp(154) := LDI & "00" & '0' & x"09";	-- LDI $9 	#Carrega o acumulador com  valor 9
tmp(155) := STA & "00" & '0' & x"0C";	-- STA @12 	#Armazena o valor das dezenas
tmp(156) := LDA & "00" & '0' & x"0D";	-- LDA @13 	#Lê o valor das centenas
tmp(157) := CEQ & "00" & '0' & x"00";	-- CEQ @0 	#Verifica se o valor das centenas é igual a 0
tmp(158) := JEQ & "00" & '0' & x"A3";	-- JEQ @163	#Se sim, decremente a unidade de milhar
tmp(159) := LDA & "00" & '0' & x"0D";	-- LDA @13 	#Carrega o acumulador com  valor 1
tmp(160) := SUB & "00" & '0' & x"01";	-- SUB @1 	#Subtrai o valor das centenas com 1
tmp(161) := STA & "00" & '0' & x"0D";	-- STA @13 	#Armazena o valor das centenas
tmp(162) := RET & "00" & '0' & x"00";	-- RET 	#Retorna ao loop principal
tmp(163) := LDI & "00" & '0' & x"09";	-- LDI $9 	#Carrega o acumulador com  valor 9
tmp(164) := STA & "00" & '0' & x"0D";	-- STA @13 	#Armazena o valor das centenas
tmp(165) := LDA & "00" & '0' & x"0E";	-- LDA @14 	#Lê o valor das unidades de milhar
tmp(166) := CEQ & "00" & '0' & x"00";	-- CEQ @0 	#Verifica se o valor das unidades de milhar é igual a 0
tmp(167) := JEQ & "00" & '0' & x"AC";	-- JEQ @172	#Se sim, decremente a dezena de milhar
tmp(168) := LDA & "00" & '0' & x"0E";	-- LDA @14 	#Carrega o acumulador com  valor 1
tmp(169) := SUB & "00" & '0' & x"01";	-- SUB @1 	#Subtrai o valor das unidades de milhar com 1
tmp(170) := STA & "00" & '0' & x"0E";	-- STA @14 	#Armazena o valor das unidades de milhar
tmp(171) := RET & "00" & '0' & x"00";	-- RET 	#Retorna ao loop principal
tmp(172) := LDI & "00" & '0' & x"09";	-- LDI $9 	#Carrega o acumulador com  valor 9
tmp(173) := STA & "00" & '0' & x"0E";	-- STA @14 	#Armazena o valor das unidades de milhar
tmp(174) := LDA & "00" & '0' & x"0F";	-- LDA @15 	#Lê o valor das dezenas de milhar
tmp(175) := CEQ & "00" & '0' & x"00";	-- CEQ @0 	#Verifica se o valor das dezenas de milhar é igual a 0
tmp(176) := JEQ & "00" & '0' & x"B5";	-- JEQ @181	#Se sim, decremente a centena de milhar
tmp(177) := LDA & "00" & '0' & x"0F";	-- LDA @15 	#Carrega o acumulador com  valor 1
tmp(178) := SUB & "00" & '0' & x"01";	-- SUB @1 	#Subtrai o valor das dezenas de milhar com 1
tmp(179) := STA & "00" & '0' & x"0F";	-- STA @15 	#Armazena o valor das dezenas de milhar
tmp(180) := RET & "00" & '0' & x"00";	-- RET 	#Retorna ao loop principal
tmp(181) := LDI & "00" & '0' & x"09";	-- LDI $9 	#Carrega o acumulador com  valor 9
tmp(182) := STA & "00" & '0' & x"0F";	-- STA @15 	#Armazena o valor das dezenas de milhar
tmp(183) := LDA & "00" & '0' & x"10";	-- LDA @16 	#Lê o valor das centenas de milhar
tmp(184) := CEQ & "00" & '0' & x"00";	-- CEQ @0 	#Verifica se o valor das centenas de milhar é igual a 0
tmp(185) := JEQ & "00" & '0' & x"BE";	-- JEQ @190	#Se sim, deixe tudo zero
tmp(186) := LDA & "00" & '0' & x"10";	-- LDA @16 	#Carrega o acumulador com  valor 1
tmp(187) := SUB & "00" & '0' & x"01";	-- SUB @1 	#Subtrai o valor das centenas de milhar com 1
tmp(188) := STA & "00" & '0' & x"10";	-- STA @16 	#Armazena o valor das centenas de milhar
tmp(189) := RET & "00" & '0' & x"00";	-- RET 	#Retorna ao loop principal
tmp(190) := LDI & "00" & '0' & x"00";	-- LDI $0 	#Carrega o acumulador com  valor 0
tmp(191) := STA & "00" & '0' & x"0B";	-- STA @11 	#Armazena o valor das unidades
tmp(192) := STA & "00" & '0' & x"0C";	-- STA @12 	#Armazena o valor das dezenas
tmp(193) := STA & "00" & '0' & x"0D";	-- STA @13 	#Armazena o valor das centenas
tmp(194) := STA & "00" & '0' & x"0E";	-- STA @14 	#Armazena o valor das unidades de milhar
tmp(195) := STA & "00" & '0' & x"0F";	-- STA @15 	#Armazena o valor das dezenas de milhar
tmp(196) := STA & "00" & '0' & x"10";	-- STA @16 	#Armazena o valor das centenas de milhar
tmp(197) := RET & "00" & '0' & x"00";	-- RET 	#Retorna ao loop principal
tmp(198) := LDA & "00" & '0' & x"0B";	-- LDA @11 	#Lê o valor das unidades
tmp(199) := STA & "00" & '1' & x"20";	-- STA @288 	#Escreve o valor das unidades em HEX0
tmp(200) := LDA & "00" & '0' & x"0C";	-- LDA @12 	#Lê o valor das dezenas
tmp(201) := STA & "00" & '1' & x"21";	-- STA @289 	#Escreve o valor das dezenas em HEX1
tmp(202) := LDA & "00" & '0' & x"0D";	-- LDA @13 	#Lê o valor das centenas
tmp(203) := STA & "00" & '1' & x"22";	-- STA @290 	#Escreve o valor das centenas em HEX2
tmp(204) := LDA & "00" & '0' & x"0E";	-- LDA @14 	#Lê o valor das unidades de milhar
tmp(205) := STA & "00" & '1' & x"23";	-- STA @291 	#Escreve o valor das unidades de milhar em HEX3
tmp(206) := LDA & "00" & '0' & x"0F";	-- LDA @15 	#Lê o valor das dezenas de milhar
tmp(207) := STA & "00" & '1' & x"24";	-- STA @292 	#Escreve o valor das dezenas de milhar em HEX4
tmp(208) := LDA & "00" & '0' & x"10";	-- LDA @16 	#Lê o valor das centenas de milhar
tmp(209) := STA & "00" & '1' & x"25";	-- STA @293 	#Escreve o valor das centenas de milhar em HEX5
tmp(210) := RET & "00" & '0' & x"00";	-- RET 	#Retorna ao loop principal
tmp(211) := STA & "00" & '1' & x"FE";	-- STA @KEY1 	#Limpa a leitura de KEY1
tmp(212) := JSR & "00" & '1' & x"11";	-- JSR @273	#Limpa os LEDs
tmp(213) := LDI & "00" & '0' & x"01";	-- LDI $1 	#Carrega o acumulador com  valor 1
tmp(214) := STA & "00" & '1' & x"00";	-- STA @256 	#Acende o LEDR0 para indicar que está configurando as unidades de segundos
tmp(215) := LDA & "00" & '1' & x"40";	-- LDA @320 	#Lê SW0-SW7
tmp(216) := STA & "00" & '1' & x"20";	-- STA @288 	#Escreve o valor das unidades de segundos em HEX0
tmp(217) := JSR & "00" & '1' & x"16";	-- JSR @278	#Chama a subrotina de comparação de KEY1
tmp(218) := JEQ & "00" & '0' & x"D7";	-- JEQ @215	#Se não foi, continue aguardando
tmp(219) := LDA & "00" & '1' & x"40";	-- LDA @320
tmp(220) := AND1 & "00" & '0' & x"2D";	-- AND1 @45
tmp(221) := STA & "00" & '0' & x"0B";	-- STA @11 	#Armazena o valor das unidades de segundos
tmp(222) := JSR & "00" & '1' & x"11";	-- JSR @273	#Limpa os LEDs
tmp(223) := STA & "00" & '1' & x"FE";	-- STA @KEY1 	#Limpa a leitura de KEY1
tmp(224) := RET & "00" & '0' & x"00";	-- RET 	#Retorna ao loop principal
tmp(225) := LDA & "00" & '0' & x"0B";	-- LDA @11 	#Lê o valor das unidades
tmp(226) := CEQ & "00" & '0' & x"15";	-- CEQ @21 	#Compara com o valor das unidades do limite
tmp(227) := JEQ & "00" & '0' & x"E5";	-- JEQ @229	#Se for igual, verifica as dezenas
tmp(228) := RET & "00" & '0' & x"00";	-- RET 	#Se for diferente, retorna ao loop principal
tmp(229) := LDA & "00" & '0' & x"0C";	-- LDA @12 	#Lê o valor das dezenas
tmp(230) := CEQ & "00" & '0' & x"16";	-- CEQ @22 	#Compara com o valor das dezenas do limite
tmp(231) := JEQ & "00" & '0' & x"E9";	-- JEQ @233	#Se for igual, verifica as centenas
tmp(232) := RET & "00" & '0' & x"00";	-- RET 	#Se for diferente, retorna ao loop principal
tmp(233) := LDA & "00" & '0' & x"0D";	-- LDA @13 	#Lê o valor das centenas
tmp(234) := CEQ & "00" & '0' & x"17";	-- CEQ @23 	#Compara com o valor das centenas do limite
tmp(235) := JEQ & "00" & '0' & x"ED";	-- JEQ @237	#Se for igual, verifica as unidades de milhar
tmp(236) := RET & "00" & '0' & x"00";	-- RET 	#Se for diferente, retorna ao loop principal
tmp(237) := LDA & "00" & '0' & x"0E";	-- LDA @14 	#Lê o valor das unidades de milhar
tmp(238) := CEQ & "00" & '0' & x"18";	-- CEQ @24 	#Compara com o valor das unidades de milhar do limite
tmp(239) := JEQ & "00" & '0' & x"F1";	-- JEQ @241	#Se for igual, verifica as dezenas de milhar
tmp(240) := RET & "00" & '0' & x"00";	-- RET 	#Se for diferente, retorna ao loop principal
tmp(241) := LDA & "00" & '0' & x"0F";	-- LDA @15 	#Lê o valor das dezenas de milhar
tmp(242) := CEQ & "00" & '0' & x"19";	-- CEQ @25 	#Compara com o valor das dezenas de milhar do limite
tmp(243) := JEQ & "00" & '0' & x"F5";	-- JEQ @245	#Se for igual, verifica as centenas de milhar
tmp(244) := RET & "00" & '0' & x"00";	-- RET 	#Se for diferente, retorna ao loop principal
tmp(245) := LDA & "00" & '0' & x"10";	-- LDA @16 	#Lê o valor das centenas de milhar
tmp(246) := CEQ & "00" & '0' & x"1A";	-- CEQ @26 	#Compara com o valor das centenas de milhar do limite
tmp(247) := JEQ & "00" & '0' & x"F9";	-- JEQ @249	#Se for igual, ative a flag de inibir contagem e ascenda o LED de limite atingido
tmp(248) := RET & "00" & '0' & x"00";	-- RET 	#Se for diferente, retorna ao loop principal
tmp(249) := LDI & "00" & '0' & x"01";	-- LDI $1 	#Carrega o acumulador com  valor 1
tmp(250) := STA & "00" & '0' & x"11";	-- STA @17 	#Ativa a flag de inibir contagem
tmp(251) := STA & "00" & '1' & x"01";	-- STA @257 	#Acende o LED de limite atingido
tmp(252) := RET & "00" & '0' & x"00";	-- RET 	#Retorna ao loop principal
tmp(253) := STA & "00" & '1' & x"FC";	-- STA @FPGA_RESET 	#Limpa a leitura de FPGA_RESET
tmp(254) := LDI & "00" & '0' & x"00";	-- LDI $0 	#Carrega o acumulador com  valor 0
tmp(255) := STA & "00" & '0' & x"0B";	-- STA @11 	#Zera o valor das unidades
tmp(256) := STA & "00" & '0' & x"0C";	-- STA @12 	#Zera o valor das dezenas
tmp(257) := STA & "00" & '0' & x"0D";	-- STA @13 	#Zera o valor das centenas
tmp(258) := STA & "00" & '0' & x"0E";	-- STA @14 	#Zera o valor das unidades de milhar
tmp(259) := STA & "00" & '0' & x"0F";	-- STA @15 	#Zera o valor das dezenas de milhar
tmp(260) := STA & "00" & '0' & x"10";	-- STA @16 	#Zera o valor das centenas de milhar
tmp(261) := STA & "00" & '0' & x"11";	-- STA @17 	#Zera a flag de inibir contagem
tmp(262) := STA & "00" & '1' & x"02";	-- STA @258 	#Apaga o LED de overflow
tmp(263) := STA & "00" & '1' & x"01";	-- STA @257 	#Apaga o LED de limite atingido
tmp(264) := RET & "00" & '0' & x"00";	-- RET 	#Retorna ao loop principal
tmp(265) := LDI & "00" & '0' & x"00";	-- LDI $0 	#Carrega o acumulador com  valor 0
tmp(266) := STA & "00" & '1' & x"20";	-- STA @288 	#Zera HEX0
tmp(267) := STA & "00" & '1' & x"21";	-- STA @289 	#Zera HEX1
tmp(268) := STA & "00" & '1' & x"22";	-- STA @290 	#Zera HEX2
tmp(269) := STA & "00" & '1' & x"23";	-- STA @291 	#Zera HEX3
tmp(270) := STA & "00" & '1' & x"24";	-- STA @292 	#Zera HEX4
tmp(271) := STA & "00" & '1' & x"25";	-- STA @293 	#Zera HEX5
tmp(272) := RET & "00" & '0' & x"00";	-- RET 	#Retorna
tmp(273) := LDI & "00" & '0' & x"00";	-- LDI $0 	#Carrega o acumulador com  valor 0
tmp(274) := STA & "00" & '1' & x"00";	-- STA @256 	#Zera dos LDR0-LDR7
tmp(275) := STA & "00" & '1' & x"01";	-- STA @257 	#Zera dos LDR8
tmp(276) := STA & "00" & '1' & x"02";	-- STA @258 	#Zera dos LDR9
tmp(277) := RET & "00" & '0' & x"00";	-- RET 	#Retorna
tmp(278) := LDA & "10" & '1' & x"61";	-- LDA R2, 353 	#Lê KEY1
tmp(279) := AND1 & "10" & '0' & x"01";	-- AND1 R2, 1 	#Mask
tmp(280) := CEQ & "10" & '0' & x"00";	-- CEQ R2, 0 	#Verifica se KEY1 não foi pressionado
tmp(281) := RET & "00" & '0' & x"00";	-- RET 	#Se Retorna




		  return tmp;
    end initMemory;

    signal memROM : blocoMemoria := initMemory;

begin
    Dado <= memROM (to_integer(unsigned(Endereco)));
end architecture;